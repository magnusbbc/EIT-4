LIBRARY IEEE; 
USE IEEE.STD_LOGIC_1164.ALL; 
USE IEEE.NUMERIC_STD.ALL; 
  
ENTITY ALU_TB IS 
END ALU_TB; 
   
ARCHITECTURE Behavioral OF ALU_TB IS 
    
  signal   operand_a    :  std_logic_vector(15 DOWNTO 0); -- Operands 1 and 2 
  signal   operand_b    :  std_logic_vector(15 DOWNTO 0); -- Operands 1 and 2   
  signal   Operation   :  std_logic_vector(5 DOWNTO 0); 
  
  signal Overflow_Flag      :  std_logic; -- Flag raised when overflow is present 
  signal Signed_Flag        :  std_logic; -- Flag that does something? 
  signal Zero_Flag          :  std_logic; -- Flag raised when operands are equal? 
  signal Parity_Flag        :  std_logic; -- Flag raised when a carry is present after adding 
  signal Carry_Flag         :  std_logic; -- Flag raised when operands are carry 
--    signal flags          :  std_logic_vector(4 downto 0); 
    signal Result             :  std_logic_vector(15 DOWNTO 0); 
     
     
  --Clock Constants 
  constant TbPeriod : time := 10 ns; 
  signal TbClock : std_logic := '0'; 
  signal TbSimEnded : std_logic := '0'; 
  signal cnt : integer := 0; 
  
BEGIN 
  ALU : ENTITY work.ALU(Behavioral)  
  PORT MAP( 
  operand_a => operand_a, 
  operand_b => operand_b, 
  operation => operation, 
  parity_Flag => parity_Flag, 
  signed_Flag => signed_Flag, 
  overflow_Flag => overflow_Flag, 
  zero_Flag => zero_Flag, 
  Carry_Flag => Carry_Flag, 
  result => result 
--  flags => flags 
  ); 
   
  -- Clock generation 
TbClock <= not TbClock after TbPeriod/2 when TbSimEnded /= '1' else '0'; 
   
stim_proc:process(TbClock) 
begin 
     
    IF(rising_edge(TbClock)) THEN 
        CASE cnt is  
            when 1 => 
              operation <= "000010";  -- Add 
              operand_a <= x"0000"; 
              operand_b <= x"0000"; 
              cnt<= cnt+1;           
            when 2 => 
              operand_a <= x"0000"; 
              operand_b <= x"2000"; 
              cnt<= cnt+1;           
            when 3 => 
              operand_a <= x"f000"; 
              operand_b <= x"1000"; 
              cnt<= cnt+1;           
            when 4 => 
              operand_a <= x"7000"; 
              operand_b <= x"5000"; 
              cnt<= cnt+1;           
            when 5 => 
              operand_a <= x"e000"; 
              operand_b <= x"b000"; 
              cnt<= cnt+1;           
            when 6 => 
              operand_a <= x"f000"; 
              operand_b <= x"f000"; 
              cnt<= cnt+1; 
            when 7 => 
              operand_a <= x"f000"; 
              operand_b <= x"8000"; 
              cnt<= cnt+1; 
            when 8 => 
              operation <= "000101"; -- AND 
              operand_a <= x"0000"; 
              operand_b <= x"0000"; 
              cnt<= cnt+1;           
            when 9 => 
              operand_a <= x"0000"; 
              operand_b <= x"5000"; 
              cnt<= cnt+1; 
            when 10 => 
              operand_a <= x"0000"; 
              operand_b <= x"A000"; 
              cnt<= cnt+1; 
            when 11 => 
              operand_a <= x"0000"; 
              operand_b <= x"FFFF"; 
              cnt<= cnt+1; 
            when 12 => 
              operand_a <= x"F000"; 
              operand_b <= x"F000"; 
              cnt<= cnt+1; 
            when 13 => 
              operation <= "000110"; -- OR 
              operand_a <= x"0000"; 
              operand_b <= x"0000"; 
              cnt<= cnt+1;           
            when 14 => 
              operand_a <= x"0000"; 
              operand_b <= x"5000"; 
              cnt<= cnt+1; 
            when 15 => 
              operand_a <= x"0000"; 
              operand_b <= x"A000"; 
              cnt<= cnt+1; 
            when 16 => 
              operand_a <= x"0000"; 
              operand_b <= x"FFFF"; 
              cnt<= cnt+1; 
            when 17 => 
              operand_a <= x"F000"; 
              operand_b <= x"F000"; 
              cnt<= cnt+1; 
            when 18 => 
              operation <= "000111"; -- XOR 
              operand_a <= x"0000"; 
              operand_b <= x"0000"; 
              cnt<= cnt+1;           
            when 19 => 
              operand_a <= x"0000"; 
              operand_b <= x"5000"; 
              cnt<= cnt+1; 
            when 20 => 
              operand_a <= x"0000"; 
              operand_b <= x"A000"; 
              cnt<= cnt+1; 
            when 21 => 
              operand_a <= x"0000"; 
              operand_b <= x"FFFF"; 
              cnt<= cnt+1; 
            when 22 => 
              operand_a <= x"F000"; 
              operand_b <= x"F000"; 
              cnt<= cnt+1; 
            when 23 => 
              operation <= "001000"; -- Negate A 
              operand_a <= x"0000"; 
              operand_b <= x"0000"; 
              cnt<= cnt+1;           
            when 24 => 
              operand_a <= x"1000"; 
              operand_b <= x"0000"; 
              cnt<= cnt+1; 
            when 25 => 
              operand_a <= x"8000"; 
              operand_b <= x"0000"; 
              cnt<= cnt+1; 
            when 26 => 
              operand_a <= x"9000"; 
              operand_b <= x"0000"; 
              cnt<= cnt+1; 
            when 27 => 
              operand_a <= x"F000"; 
              operand_b <= x"0000"; 
              cnt<= cnt+1; 
            when 28 => 
               operand_a <= x"0000"; 
               operand_b <= x"F000"; 
               cnt<= cnt+1;           
            when 29 => 
               operand_a <= x"1000"; 
               operand_b <= x"F000"; 
               cnt<= cnt+1; 
            when 30 => 
               operand_a <= x"8000"; 
               operand_b <= x"F000"; 
               cnt<= cnt+1; 
            when 31 => 
               operand_a <= x"9000"; 
               operand_b <= x"F000"; 
               cnt<= cnt+1; 
            when 32 => 
               operand_a <= x"F000"; 
               operand_b <= x"F000"; 
               cnt<= cnt+1; 
            when 33 => 
               operation <= "001001"; -- Negate B 
               operand_b <= x"0000"; 
               operand_a <= x"0000"; 
               cnt<= cnt+1;           
            when 34 => 
               operand_b <= x"1000"; 
               operand_a <= x"0000"; 
               cnt<= cnt+1; 
            when 35 => 
               operand_b <= x"8000"; 
               operand_a <= x"0000"; 
               cnt<= cnt+1; 
            when 36 => 
               operand_b <= x"9000"; 
               operand_a <= x"0000"; 
               cnt<= cnt+1; 
            when 37 => 
               operand_b <= x"F000"; 
               operand_a <= x"0000"; 
               cnt<= cnt+1; 
            when 38 => 
                operand_b <= x"0000"; 
                operand_a <= x"F000"; 
                cnt<= cnt+1;           
            when 39 => 
                operand_b <= x"1000"; 
                operand_a <= x"F000"; 
                cnt<= cnt+1; 
            when 40 => 
                operand_b <= x"8000"; 
                operand_a <= x"F000"; 
                cnt<= cnt+1; 
            when 41 => 
                operand_b <= x"9000"; 
                operand_a <= x"F000"; 
                cnt<= cnt+1; 
            when 42 => 
                operand_b <= x"F000"; 
                operand_a <= x"F000"; 
                cnt<= cnt+1; 
            when 43 => 
                operation <= "001010"; -- NOT A 
                operand_a <= x"0000"; 
                operand_b <= x"0000"; 
                cnt<= cnt+1;           
            when 44 => 
                operand_a <= x"5000"; 
                operand_b <= x"0000"; 
                cnt<= cnt+1; 
            when 45 => 
                operand_a <= x"A000"; 
                operand_b <= x"0000"; 
                cnt<= cnt+1; 
            when 46 => 
                operand_a <= x"FFFF"; 
                operand_b <= x"0000"; 
                cnt<= cnt+1; 
            when 47 => 
                operand_a <= x"0000"; 
                operand_b <= x"F000"; 
                cnt<= cnt+1; 
            when 48 => 
                operand_a <= x"5000"; 
                operand_b <= x"F000"; 
                cnt<= cnt+1;           
            when 49 => 
                operand_a <= x"A000"; 
                operand_b <= x"F000"; 
                cnt<= cnt+1; 
            when 50 => 
                operand_a <= x"FFFF"; 
                operand_b <= x"F000"; 
                cnt<= cnt+1; 
            when 51 => 
                operation <= "001011"; -- NOT B             
                operand_a <= x"0000"; 
                operand_b <= x"0000"; 
                cnt<= cnt+1; 
            when 52 => 
                operand_a <= x"0000"; 
                operand_b <= x"5000"; 
                cnt<= cnt+1; 
            when 53 => 
                operand_a <= x"0000"; 
                operand_b <= x"A000"; 
                cnt<= cnt+1;           
            when 54 => 
                operand_a <= x"0000"; 
                operand_b <= x"FFFF"; 
                cnt<= cnt+1; 
            when 55 => 
                operand_a <= x"F000"; 
                operand_b <= x"0000"; 
                cnt<= cnt+1; 
            when 56 => 
                operand_a <= x"F000"; 
                operand_b <= x"5000"; 
                cnt<= cnt+1; 
            when 57 => 
                operand_a <= x"F000"; 
                operand_b <= x"A000"; 
                cnt<= cnt+1; 
            when 58 => 
                operand_a <= x"F000"; 
                operand_b <= x"FFFF"; 
                 cnt<= cnt+1;           
            when 59 => 
                operation <= "001100"; -- Logic left shift  
                operand_a <= x"0000"; 
                operand_b <= x"0000"; 
                 cnt<= cnt+1; 
            when 60 => 
                operand_a <= x"0001"; 
                operand_b <= x"0000"; 
                 cnt<= cnt+1; 
            when 61 => 
                operand_a <= x"0001"; 
                operand_b <= x"0001"; 
                 cnt<= cnt+1; 
            when 62 => 
                operand_a <= x"0001"; 
                operand_b <= x"000F"; 
                 cnt<= cnt+1; 
            when 63 => 
                operand_a <= x"0001"; 
                operand_b <= x"0010"; 
                 cnt<= cnt+1;           
            when 64 => 
                operation <= "001101"; -- Logic right shift  
                operand_a <= x"0000"; 
                operand_b <= x"0000"; 
                 cnt<= cnt+1; 
            when 65 => 
                operand_a <= x"8000"; 
                operand_b <= x"0000"; 
                 cnt<= cnt+1; 
            when 66 => 
                operand_a <= x"8000"; 
                operand_b <= x"0001"; 
                 cnt<= cnt+1; 
            when 67 => 
                operand_a <= x"8000"; 
                operand_b <= x"000F"; 
                 cnt<= cnt+1; 
            when 68 => 
                operand_a <= x"8000"; 
                operand_b <= x"0010"; 
                  cnt<= cnt+1;           
            when 69 => 
                operation <= "001110"; -- Arith right shift  
                operand_a <= x"0000"; 
                operand_b <= x"0000"; 
                  cnt<= cnt+1; 
            when 70 => 
                operand_a <= x"8000"; 
                operand_b <= x"0000"; 
                  cnt<= cnt+1; 
            when 71 => 
                operand_a <= x"8000"; 
                operand_b <= x"0001"; 
                  cnt<= cnt+1; 
            when 72 => 
                operand_a <= x"8000"; 
                operand_b <= x"000F"; 
                  cnt<= cnt+1; 
            when 73 => 
                operand_a <= x"8000"; 
                operand_b <= x"0010"; 
                  cnt<= cnt+1;           
            when 74 => 
                operand_a <= x"4000"; 
                operand_b <= x"0001"; 
                  cnt<= cnt+1; 
            when 75 => 
                operand_a <= x"4000"; 
                operand_b <= x"000E"; 
                  cnt<= cnt+1; 
            when 76 => 
                operand_a <= x"4000"; 
                operand_b <= x"000F"; 
                  cnt<= cnt+1; 
            when 77 => 
                operation <= "001111"; -- Pass A 
                operand_a <= x"0000"; 
                operand_b <= x"0000"; 
                  cnt<= cnt+1; 
            when 78 => 
                operand_a <= x"5000"; 
                operand_b <= x"0000"; 
                   cnt<= cnt+1;           
            when 79 => 
                operand_a <= x"FFFF"; 
                operand_b <= x"0000"; 
                   cnt<= cnt+1; 
            when 80 => 
                operand_a <= x"0000"; 
                operand_b <= x"F000"; 
                cnt<= cnt+1; 
            when 81 => 
                operand_a <= x"5000"; 
                operand_b <= x"F000"; 
                cnt<= cnt+1; 
            when 82 => 
                operand_a <= x"FFFF"; 
                operand_b <= x"F000"; 
                cnt<= cnt+1; 
            when 83 => 
                operation <= "010000"; -- Pass B  
                operand_a <= x"0000"; 
                operand_b <= x"0000"; 
                cnt<= cnt+1; 
            when 84 => 
                operand_a <= x"0000"; 
                operand_b <= x"5000"; 
                cnt<= cnt+1; 
            when 85 => 
                operand_a <= x"0000"; 
                operand_b <= x"F000"; 
                   cnt<= cnt+1;           
            when 86 => 
                operand_a <= x"F000"; 
                operand_b <= x"0000"; 
                   cnt<= cnt+1; 
            when 87 => 
                operand_a <= x"F000"; 
                operand_b <= x"5000"; 
                cnt<= cnt+1; 
            when 88 => 
                operand_a <= x"F000"; 
                operand_b <= x"F000"; 
                cnt<= cnt+1; 
            when 89 => 
                operation <= "010001"; -- INC A  
                operand_a <= x"0000"; 
                operand_b <= x"0000"; 
                   cnt<= cnt+1; 
            when 90 => 
                operand_a <= x"FFFF"; 
                operand_b <= x"0000"; 
                   cnt<= cnt+1; 
            when 91 => 
                operand_a <= x"4000"; 
                operand_b <= x"0000"; 
                   cnt<= cnt+1; 
            when 92 => 
                operation <= "010010"; --INC B 
                operand_a <= x"0000"; 
                operand_b <= x"0000"; 
                   cnt<= cnt+1;           
            when 93 => 
                operand_a <= x"0000"; 
                operand_b <= x"FFFF"; 
                   cnt<= cnt+1; 
            when 94 => 
                operand_a <= x"0000"; 
                operand_b <= x"4000"; 
                   cnt<= cnt+1; 
            when 95 => 
                operation <= "010011"; --NOP 
                operand_a <= x"0000"; 
                operand_b <= x"F000"; 
                   cnt<= cnt+1;  
            when 96 => 
                operation <= "000011"; --SUB 
                operand_a <= x"0000"; 
                operand_b <= x"0000"; 
                   cnt<= cnt+1; 
            when 97 => 
                operand_a <= x"0014"; 
                operand_b <= x"000A"; 
                cnt<= cnt+1; 
            when 98 => 
                operand_a <= x"000A"; 
                operand_b <= x"0014"; 
                cnt<= cnt+1; 
            when 99 => 
                operand_a <= x"FFF6"; 
                operand_b <= x"0014"; 
                   cnt<= cnt+1; 
            when 100 => 
                operand_a <= x"FFF6"; 
                operand_b <= x"FFEC"; 
                   cnt<= cnt+1; 
            when 101 => 
                operand_a <= x"FFEC"; 
                operand_b <= x"FFF6"; 
                   cnt<= cnt+1; 
            when 102 => 
                operand_a <= x"8000"; 
                operand_b <= x"7000"; 
                   cnt<= cnt+1;           
            when 103 => 
                operation <= "000100";  --MULT 
                operand_a <= x"0000"; 
                operand_b <= x"0000"; 
                   cnt<= cnt+1; 
            when 104 => 
                operand_a <= x"7000"; 
                operand_b <= x"0001"; 
                   cnt<= cnt+1; 
            when 105 => 
                operand_a <= x"FFFE"; 
                operand_b <= x"0002"; 
                   cnt<= cnt+1;  
            when 106 => 
                operand_a <= x"7000"; 
                operand_b <= x"0005"; 
                   cnt<= cnt+1; 
            when 107 => 
                operand_a <= x"E000"; 
                operand_b <= x"FFFE"; 
                   cnt<= cnt+1;           
            when 108 => 
                operand_a <= x"C000"; 
                operand_b <= x"FFFA"; 
                   cnt<= cnt+1; 
                            
            when others =>  
              cnt<= cnt+1; 
        End case;      
        IF(cnt = 108) THEN 
            TbSimEnded <= '1'; 
            --wait; 
        END IF;  
    END IF; 
end process; 
  
   
END Behavioral;