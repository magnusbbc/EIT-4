#include "Config.hvhd"
--------------------------------------------------------------------------------------
--Engineer: Magnus Christensen
--Module Name: Master
--
--Description:
--
--
--
--------------------------------------------------------------------------------------


--Definition of control lines
#define ALU_CONTROL 18 DOWNTO 13
#define JUMP_CONTROL 12 DOWNTO 10
#define MEMORY_READ 9
#define MEMORY_WRITE 8
#define REGISTER_WRITE 7
#define MEMORY_WRITE_BACK 6
#define IMMEDIATE_SELECT 5
#define PUSH 4
#define POP 3
#define SWITCH_READ_WRITE 2
#define MEMORY_TO_PC 1
#define HALT 0

--definition of instruction lines
#define OPCODE 31 DOWNTO 26
#define REGISTER_READ_INDEX_1 25 DOWNTO 21
#define REGISTER_READ_INDEX_2 15 DOWNTO 11
#define REGISTER_WRITE_INDEX_1 20 DOWNTO 16
#define IMMEDIATE 15 DOWNTO 0

#define PUSH_PC "10000100000000001111100000000000"
#define POP_PC "10000000000111110000000000000000"

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_unsigned.ALL;
USE IEEE.NUMERIC_STD.ALL;


ENTITY Master IS
	PORT (
		clk : IN std_logic;
		btn : IN std_logic_vector(2 DOWNTO 0);
		sseg : OUT std_logic_vector(31 DOWNTO 0);
		led : OUT std_logic_vector(9 DOWNTO 0);
		
		bclk   : IN std_logic := '0';
		ws     : IN std_logic := '0';
		Din    : IN std_logic := '0';
		
		bclkO     : out std_logic := '0';
		wsO       : out std_logic := '0';
		DOut : out std_logic := '0'
	);
END ENTITY Master;

ARCHITECTURE Behavioral OF Master IS
	SIGNAL btn_inverted : std_logic_vector(2 DOWNTO 0) := "000";
	--Control and instruction registers
	SIGNAL control_signals : Std_logic_vector(CONTROL_SIZE DOWNTO 0); --Control signals generated by the control block
	SIGNAL instruction : std_logic_vector(INSTRUCTION_SIZE DOWNTO 0); --Instruction sent to the system
	SIGNAL pram_data_out : std_logic_vector(INSTRUCTION_SIZE DOWNTO 0); --Instruction outputted by the program memory
	
	--Wires
	SIGNAL operand_a, operand_b, alu_output : std_logic_vector(WORD_SIZE DOWNTO 0); -- ALU inputs and output wires
	SIGNAL stack_controller_out : std_logic_vector(WORD_SIZE DOWNTO 0); --Stackpointer address wires
	SIGNAL register_writeback : std_logic_vector(WORD_SIZE DOWNTO 0); --Wires to connect ALU/Memory output to register writeback logic
	SIGNAL dram_address_index : std_logic_vector(WORD_SIZE DOWNTO 0); --Wires connected to the memory controllers address port
	SIGNAL r2_w1_switch : std_logic_vector(4 DOWNTO 0); --Size '5' to be able to index register. Is used to switch between indexing Read_2 and Write_1 register

	--PRAM Signals
	SIGNAL pc : std_logic_vector(9 DOWNTO 0) := (OTHERS => '0'); --Program Counter
	SIGNAL pram_address_index : std_logic_vector(9 DOWNTO 0) := (OTHERS => '0'); --Wires connected to the PRAM's address port
	SIGNAL pc_alt : std_logic_vector(9 DOWNTO 0) := (OTHERS => '0'); --Alternative new PC (e.g. ALU/Memory Output), used when changing the PC (for jumps)
	SIGNAL interrupt_address : std_logic_vector(9 DOWNTO 0) := (OTHERS => '0'); --Interrupt address, address that the ISR points to
	SIGNAL pram_data_in : std_logic_vector(INSTRUCTION_SIZE DOWNTO 0); --Not used in current implementation, used to write to program memory
	SIGNAL pram_write_enable : std_logic := '0'; --Program memory write enable disabled in current implementation
	SIGNAL pram_read_enable : std_logic := '1'; --Program memory read enable always on in current implementation
	--DRAM Signals
	SIGNAL dram_data_out : std_logic_vector(WORD_SIZE DOWNTO 0); --Data RAM output data
	SIGNAL dram_data_in : std_logic_vector(WORD_SIZE DOWNTO 0); --Data RAM Input data, either source_register_2_output, or --- (needed for proper interrupt implementation)

	--Reg Signals
	SIGNAL source_register_2_output : STD_logic_vector(WORD_SIZE DOWNTO 0); --2nd indexed register output, needed as a buffer to be able to switch bewtween register_2 and Immediate input to the alu

	SIGNAL jmp_enable : std_logic := '0'; --Is '0' when PC increments by 1, is set to '1' when jump occours
	SIGNAL pc_overwrite, sp_overwrite : std_logic := '0'; --SP and PC are special registers, and PC/sp_overwrite needs to be '1' to be able to change their values

	SIGNAL pc_register_file_input : std_logic_vector(WORD_SIZE DOWNTO 0); --Routes PC+1 into the register file

	SIGNAL interrupt_cpu : std_logic := '0'; --Interrupt signal for the CPU
	SIGNAL Interrupt_latch : std_logic := '0'; --Latch for the interrupt signal, ensures signal stays on for an additional clock cycle
	SIGNAl interrupt_enable : std_logic := '1';
	SIGNAL interrupt_nest_enable : std_logic := '1';
	SIGNAL interrupt_nest_enable_latch : std_logic := '0';

	SIGNAL pc_interrupt_push : std_logic_vector(9 DOWNTO 0) := (OTHERS => '0');
	--FLAGS
	SIGNAL parity_flag : std_logic := '0';
	SIGNAL signed_flag : std_logic := '0';
	SIGNAL overflow_flag : std_logic := '0';
	SIGNAL zero_flag : std_logic := '0';
	SIGNAL carry_flag : std_logic := '0';

	--FLAG LATCHES
	SIGNAL parity_flag_latch : std_logic := '0';
	SIGNAL signed_flag_latch : std_logic := '0';
	SIGNAL overflow_flag_latch : std_logic := '0';
	SIGNAL zero_flag_latch : std_logic := '0';
	SIGNAL carry_flag_latch : std_logic := '0';
	
	SIGNAL sys_clk : std_logic; --Clock that controls the system, can either be assigned to the normal clock (for simulation), or pll_tmp_clk
	SIGNAL pll_clk : std_logic; --PLL Clock
	SIGNAL pll_lock : std_logic; --PLL lock signal
	SIGNAL pll_tmp_clk : Std_logic; --Is assigned the pll_clk when pll_lock is detected
	SIGNAL clk_counter : std_logic_vector(24 DOWNTO 0); --Clock divider, used to switch LED (works as a clock heart beat)

BEGIN

	PLL : ENTITY work.PLL(SYN)
		PORT MAP(
			inclk0 => clk,
			c0 => pll_clk,
			locked => pll_lock
		);
	MEMCNT : ENTITY work.MemoryController
		PORT MAP(
			write_enable => control_signals(MEMORY_WRITE),
			read_enable => control_signals(MEMORY_READ),
			address => dram_address_index,
			data_in => dram_data_in,
			DO => dram_data_out,
			clk => sys_clk,
			btn => btn_inverted,
			seven_seg_control_signals => sseg,
			interrupt_address => interrupt_address,
			interrupt_cpu => interrupt_cpu,
			interrupt_enable => interrupt_enable,
			interrupt_nest_enable => interrupt_nest_enable,
			i2s_bit_clk => bclk,
			i2s_word_select => ws,
			i2s_data_in => Din,
			i2s_bit_clk_out => bclkO,
			i2s_word_select_out => wsO,
			i2s_data_out => DOut
		);

	CONTROLLER : ENTITY work.Control(Behavioral)
		PORT MAP(
			opcode => instruction(OPCODE),
			control_signals => control_signals
		);
	
	STACK : ENTITY work.Stack(Behavioral)
		PORT MAP(
			pop => control_signals(POP),
			push => control_signals(PUSH),
			clk => sys_clk,
			address_out => stack_controller_out,
			address_in => register_writeback,
			write_back => sp_overwrite
		);

	ALU : ENTITY work.ALU(Behavioral)
		PORT MAP(
			operation => control_signals(ALU_CONTROL),
			operand_a => operand_a,
			operand_b => operand_b,
			result => alu_output,
			parity_flag => parity_flag,
			signed_flag => signed_flag,
			overflow_flag => overflow_flag,
			zero_flag => zero_flag,
			carry_flag => carry_flag
		);
	PRAM : ENTITY work.MemAuto(SYN)
		PORT MAP(
			data => pram_data_in,
			q => pram_data_out,
			address => pram_address_index,
			wren => pram_write_enable,
			rden => pram_read_enable,
			clock => sys_clk
		);
	REGS : ENTITY work.RegistryInternal(Behavioral)
		PORT MAP(
			read_register_a_index => instruction(REGISTER_READ_INDEX_1),
			write_register_index => instruction(REGISTER_WRITE_INDEX_1),
			read_register_b_index => r2_w1_switch,

			register_file_data_in => register_writeback,

			register_file_data_out_a => operand_a,
			register_file_data_out_b => source_register_2_output,

			pc_value_input => pc_register_file_input,
			sp_value_input => stack_controller_out,

			write_enable => control_signals(REGISTER_WRITE),

			clk => sys_clk
		);


	WITH Interrupt_latch SELECT dram_data_in <=
	std_logic_vector(to_unsigned(to_integer(unsigned(pc_interrupt_push)),dram_data_in'length))  WHEN '1',
	source_register_2_output WHEN OTHERS;


	WITH control_signals(IMMEDIATE_SELECT) SELECT operand_b <= -- Selects Register output 2 or Immediate
	source_register_2_output WHEN '0',
	instruction(IMMEDIATE) WHEN '1',
	source_register_2_output WHEN OTHERS;

	WITH control_signals(SWITCH_READ_WRITE) SELECT r2_w1_switch <= --if SWITCH_READ_WRITE, Read 2 index will be write 1 index
	instruction(REGISTER_WRITE_INDEX_1) WHEN '1',
	instruction(REGISTER_READ_INDEX_2) WHEN OTHERS;
	
	WITH control_signals(MEMORY_WRITE_BACK) SELECT register_writeback <=
	dram_data_out WHEN '1',
	alu_output WHEN OTHERS;

	WITH to_integer(unsigned(instruction(REGISTER_WRITE_INDEX_1))) SELECT pc_overwrite <=
	'1' WHEN 31,
	'0' WHEN OTHERS;

	PROCESS (instruction(REGISTER_WRITE_INDEX_1),control_signals(SWITCH_READ_WRITE))
	BEGIN
	IF(to_integer(unsigned(instruction(REGISTER_WRITE_INDEX_1))) = 30 AND control_signals(SWITCH_READ_WRITE) /= '1') THEN
		sp_overwrite <= '1';
	ELSE
		sp_overwrite <= '0';
	END IF;
	END PROCESS;


	PROCESS(control_signals(POP),control_signals(PUSH),stack_controller_out,alu_output)
		VARIABLE TMP : std_logic_vector(1 downto 0);
	BEGIN
		TMP := control_signals(POP) & control_signals(PUSH);
		IF(to_integer(UNSIGNED(TMP)) > 0) THEN
			dram_address_index <= stack_controller_out;
		ELSE
			dram_address_index <= alu_output;
		END IF;
	END PROCESS;

	WITH to_integer(unsigned(Interrupt_latch & pc_overwrite & control_signals(JUMP_CONTROL))) SELECT jmp_enable <= --Controls branching/changing PC
	'0' WHEN 0,
	'1' WHEN 1,
	zero_flag_latch WHEN 2,
	carry_flag_latch WHEN 3,
	NOT zero_flag_latch WHEN 4,
	'1' WHEN 8, --WHEN pc_overwrite is set
	'1' WHEN 16,
	'0' WHEN OTHERS;

	PROCESS(interrupt_cpu,Interrupt_latch,control_signals(MEMORY_TO_PC),dram_data_out(9 DOWNTO 0),alu_output(9 DOWNTO 0))
	BEGIN
		IF(interrupt_cpu = '1' OR Interrupt_latch = '1') THEN
			pc_alt <= interrupt_address;
		ELSIF(control_signals(MEMORY_TO_PC) = '1') THEN
			pc_alt <= dram_data_out(9 DOWNTO 0);
		ELSE
			pc_alt <= alu_output(9 DOWNTO 0);
		END IF;
	END PROCESS;

	WITH jmp_enable SELECT pram_address_index <= --Choses instruction to be loaded based on branching
		pc_alt WHEN '1',
		pc WHEN OTHERS;



	PROCESS  (Interrupt_latch, pram_data_out)--Changes instruction if interrupt is detected
	BEGIN
		IF(Interrupt_latch = '1') THEN
			instruction <= PUSH_PC;
		ELSE
			instruction <= pram_data_out;
		END IF;
	END PROCESS;


	RUN : PROCESS (sys_clk) --Chose new value of PC based on branching
	BEGIN
		IF (rising_edge(sys_clk)) THEN --clk
			IF (Interrupt_latch = '1' AND jmp_enable /= '1') THEN
				pc <= pc;
			ELSIF (Interrupt_latch = '1' AND jmp_enable = '1') THEN
				pc <= std_logic_vector(unsigned(pc_alt) + 1);
			ELSIF (jmp_enable /= '1') THEN
				pc <= std_logic_vector(unsigned(pc) + 1);
			ELSE
				pc <= std_logic_vector(unsigned(pc_alt) + 1);
			END IF;
		END IF;
	END PROCESS;

	PROCESS(instruction, interrupt_nest_enable)
	BEGIN
		IF(interrupt_nest_enable = '0' AND interrupt_nest_enable_latch = '0') THEN
			interrupt_enable <= '0';
			interrupt_nest_enable_latch <= '1';
		ELSIF(instruction = POP_PC) THEN
			interrupt_enable <= '1';
			interrupt_nest_enable_latch <= '0';
		END IF;
	END PROCESS;

	PROCESS(sys_clk)
	BEGIN
		IF(rising_edge(sys_clk)) THEN
			IF(interrupt_cpu = '1') THEN
				Interrupt_latch <= '1';
				IF(jmp_enable = '1') THEN
					pc_interrupt_push <= std_logic_vector(unsigned(pc) - 1);
				ELSE
					pc_interrupt_push <= pc;
				END IF;
			ELSIF(Interrupt_latch = '1') THEN
				Interrupt_latch <= '0';
			END IF;
		END IF;
	END PROCESS;

	--Latches Flags in tempo register, neccesarry due to clock timing
	LATCH : PROCESS (sys_clk)
	BEGIN
		IF (rising_edge(sys_clk)) THEN
			zero_flag_latch <= zero_flag;
			overflow_flag_latch <= overflow_flag;
			signed_flag_latch <= signed_flag;
			parity_flag_latch <= parity_flag;
			carry_flag_latch <= carry_flag;
		END IF;
	END PROCESS;

	pc_register_file_input <= "000000" & std_logic_vector(unsigned(pc) + 1);

--Below controls Clock---

	WITH control_signals(HALT) SELECT sys_clk <=
	pll_tmp_clk WHEN '0',
	--DBtn(2) when '0',
	--clk when '0',
	'0' WHEN OTHERS;

	WITH pll_lock SELECT pll_tmp_clk <=
		pll_clk WHEN '1',
		'0' WHEN OTHERS;
	PROCESS (pll_clk)

	BEGIN
		IF (rising_edge(pll_clk)) THEN
			clk_counter <= std_logic_vector(unsigned(clk_counter) + 1);
		END IF;
	END PROCESS;

	btn_inverted <= not btn;

	LED(9) <= zero_flag;
	LED(8) <= overflow_flag;
	LED(7) <= signed_flag;
	LED(6) <= parity_flag;
	LED(5) <= btn_inverted(0);

	LED(0) <= clk_counter(24);
	LED(1) <= control_signals(HALT);

END ARCHITECTURE Behavioral;