-- Package Declaration Section
package Constants is
	constant ADDVAL : integer := 1;
end package Constants;