#include "Config.hvhd"

--Definition of control lines
#define ALU_CONTROL 18 DOWNTO 13
#define JUMP_CONTROL 12 DOWNTO 10
#define MEMORY_READ 9
#define MEMORY_WRITE 8
#define REGISTER_WRITE 7
#define MEMORY_WRITE_BACK 6
#define IMMEDIATE_SELECT 5
#define PUSH 4
#define POP 3
#define SWITCH_READ_WRITE 2
#define MEMORY_TO_PC 1
#define HALT 0

--definition of instruction lines
#define OPCODE 31 DOWNTO 26
#define REGISTER_READ_INDEX_1 25 DOWNTO 21
#define REGISTER_READ_INDEX_2 15 DOWNTO 11
#define REGISTER_WRITE_INDEX_1 20 DOWNTO 16
#define IMMEDIATE 15 DOWNTO 0

#define PUSH_PC "10000100000000001111100000000000"
#define POP_PC "10000000000111110000000000000000"

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_unsigned.ALL;
USE IEEE.NUMERIC_STD.ALL;


ENTITY Master IS
	PORT (
		clk : IN std_logic;
		btn : IN std_logic_vector(2 DOWNTO 0);
		sseg : OUT std_logic_vector(31 DOWNTO 0);
		led : OUT std_logic_vector(9 DOWNTO 0);
		
		bclk   : IN std_logic := '0';
		ws     : IN std_logic := '0';
		Din    : IN std_logic := '0';
		
		bclkO     : out std_logic := '0';
		wsO       : out std_logic := '0';
		DOut : out std_logic := '0'
	);
END ENTITY Master;

ARCHITECTURE Behavioral OF Master IS
	SIGNAL btn_inverted : std_logic_vector(2 DOWNTO 0) := "000";
	--Control and instruction registers
	SIGNAL CONTROL : Std_logic_vector(CONTROL_SIZE DOWNTO 0); --Control signals generated by the control block
	SIGNAL INSTRUCTION : std_logic_vector(INSTRUCTION_SIZE DOWNTO 0); --Instruction sent to the system
	SIGNAL INSTRUCTION_PRAM : std_logic_vector(INSTRUCTION_SIZE DOWNTO 0); --Instruction oututted by the program memory
	
	--Wires
	SIGNAL OP1, OP2, ALU_OUTPUT : std_logic_vector(WORD_SIZE DOWNTO 0); -- ALU inputs and output wires
	SIGNAL SP_OUT : std_logic_vector(WORD_SIZE DOWNTO 0); --Stackpointer address wires
	SIGNAL REGISTER_WRITEBACK : std_logic_vector(WORD_SIZE DOWNTO 0); --Wires to connect ALU/Memory output to register writeback logic
	SIGNAL MEM_ADDRESS : std_logic_vector(WORD_SIZE DOWNTO 0); --Wires connected to the memory controllers address port
	SIGNAL RWSWITCH : std_logic_vector(4 DOWNTO 0); --Size '5' to be able to index register. Is used to switch between indexing Read_2 and Write_1 register

	--PRAM Signals
	SIGNAL PC : std_logic_vector(9 DOWNTO 0) := (OTHERS => '0'); --Program Counter
	SIGNAL ADDR : std_logic_vector(9 DOWNTO 0) := (OTHERS => '0'); --Wires connected to the PRAM's address port
	SIGNAL PC_ALT : std_logic_vector(9 DOWNTO 0) := (OTHERS => '0'); --Alternative new PC (e.g. ALU/Memory Output), used when changing the PC (for jumps)
	SIGNAL Interrupt_addr : std_logic_vector(9 DOWNTO 0) := (OTHERS => '0'); --Interrupt address, address that the ISR points to
	SIGNAL pDataIn : std_logic_vector(INSTRUCTION_SIZE DOWNTO 0); --Not used in current implementation, used to write to program memory
	SIGNAL pDataOut : std_logic_vector(INSTRUCTION_SIZE DOWNTO 0); --Program Memory instruction output
	SIGNAL PWE : std_logic := '0'; --Program memory write enable disabled in current implementation
	SIGNAL PRE : std_logic := '1'; --Program memory read enable always on in current implementation
	--DRAM Signals
	SIGNAL dDataOut : std_logic_vector(WORD_SIZE DOWNTO 0); --Data RAM output data
	SIGNAL dDataIn : std_logic_vector(WORD_SIZE DOWNTO 0); --Data RAM Input data, either R2O, or R2O-2 (needed for proper interrupt implementation)

	--Reg Signals
	SIGNAL R2O : STD_logic_vector(WORD_SIZE DOWNTO 0); --2nd indexed register output, needed as a buffer to be able to switch bewtween register_2 and Immediate input to the alu

	SIGNAL JMP_SELECT : std_logic := '0'; --Is '0' when PC increments by 1, is set to '1' when jump occours
	SIGNAL PC_OVERWRITE, SP_OVERWRITE : std_logic := '0'; --SP and PC are special registers, and PC/SP_OVERWRITE needs to be '1' to be able to change their values

	SIGNAL PC_REG_IN : std_logic_vector(WORD_SIZE DOWNTO 0); --Routes PC+1 into the register file

	SIGNAL Interrupt_CPU : std_logic := '0'; --Interrupt signal for the CPU
	SIGNAL Interrupt_latch : std_logic := '0'; --Latch for the interrupt signal, ensures signal stays on for an additional clock cycle
	SIGNAl Interrupt_enable : std_logic := '1';
	SIGNAL Interrupt_nest_enable : std_logic := '1';
	SIGNAL Interrupt_nest_enable_latch : std_logic := '0';

	SIGNAL PC_INT_TMP : std_logic_vector(9 DOWNTO 0) := (OTHERS => '0');
	--FLAGS
	SIGNAL Parity_Flag : std_logic := '0';
	SIGNAL Signed_Flag : std_logic := '0';
	SIGNAL Overflow_Flag : std_logic := '0';
	SIGNAL Zero_Flag : std_logic := '0';
	SIGNAL Carry_Flag : std_logic := '0';

	--FLAG LATCHES
	SIGNAL Parity_Flag_Latch : std_logic := '0';
	SIGNAL Signed_Flag_Latch : std_logic := '0';
	SIGNAL Overflow_Flag_Latch : std_logic := '0';
	SIGNAL Zero_Flag_Latch : std_logic := '0';
	SIGNAL Carry_Flag_Latch : std_logic := '0';
	
	SIGNAL subClock : std_logic; --Clock that controls the system, can either be assigned to the normal clock (for simulation), or PLL_CLOCK_TEMP
	SIGNAL PLL_CLOCK : std_logic; --PLL Clock
	SIGNAL PLL_LOCK : std_logic; --PLL lock signal
	SIGNAL PLL_CLOCK_TEMP : Std_logic; --Is assigned the PLL_CLOCK when PLL_LOCK is detected
	SIGNAL DIVIDER : std_logic_vector(25 DOWNTO 0); --Clock divider, used to switch LED (works as a clock heart beat)

BEGIN

	PLL : ENTITY work.PLL(SYN)
		PORT MAP(
			inclk0 => clk,
			c0 => PLL_CLOCK,
			locked => PLL_LOCK
		);
	MEMCNT : ENTITY work.MemoryController
		PORT MAP(
			WE => CONTROL(MEMORY_WRITE),
			RE => CONTROL(MEMORY_READ),
			Address => MEM_ADDRESS,
			DI => dDataIn,
			DO => dDataOut,
			CLK => subClock,
			btn => btn_inverted,
			ss => sseg,
			control => Interrupt_addr,
			interrupt_cpu => Interrupt_CPU,
			Interrupt_enable => Interrupt_enable,
			Interrupt_nest_enable => Interrupt_nest_enable,
			bclk => bclk,
			ws => ws,
			Din => Din,
			bclkO => bclkO,
			wsO => wsO,
			DOut => DOut
		);

	CONTROLLER : ENTITY work.Control(Behavioral)
		PORT MAP(
			opcode => INSTRUCTION(OPCODE),
			cntSignal => CONTROL
		);
	
	STACK : ENTITY work.Stack(Behavioral)
		PORT MAP(
			pop => CONTROL(POP),
			push => CONTROL(PUSH),
			clk => subClock,
			addressOut => SP_OUT,
			addressIn => REGISTER_WRITEBACK,
			writeBack => SP_OVERWRITE
		);

	ALU : ENTITY work.ALU(Behavioral)
		PORT MAP(
			Operation => CONTROL(ALU_CONTROL),
			Operand1 => OP1,
			Operand2 => OP2,
			Result => ALU_OUTPUT,
			Parity_Flag => Parity_Flag,
			Signed_Flag => Signed_Flag,
			Overflow_Flag => Overflow_Flag,
			Zero_Flag => Zero_Flag,
			Carry_Flag => Carry_Flag
		);
	PRAM : ENTITY work.MemAuto(SYN)
		PORT MAP(
			data => pDataIn,
			q => INSTRUCTION_PRAM,
			address => ADDR,
			wren => PWE,
			rden => PRE,
			clock => subClock
		);
	REGS : ENTITY work.RegistryInternal(Behavioral)
		PORT MAP(
			readOne => INSTRUCTION(REGISTER_READ_INDEX_1),
			WriteOne => INSTRUCTION(REGISTER_WRITE_INDEX_1),
			readTwo => RWSWITCH,

			dataInOne => REGISTER_WRITEBACK,

			dataOutOne => OP1,
			dataOutTwo => R2O,

			pcIn => PC_REG_IN,
			spIN => SP_OUT,

			WR1_E => CONTROL(REGISTER_WRITE),

			clk => subClock
		);


	WITH Interrupt_latch SELECT dDataIn <=
	std_logic_vector(to_unsigned(to_integer(unsigned(PC_INT_TMP)),dDataIn'length))  WHEN '1',
	R2O WHEN OTHERS;


	WITH CONTROL(IMMEDIATE_SELECT) SELECT OP2 <= -- Selects Register output 2 or Immediate
	R2O WHEN '0',
	INSTRUCTION(IMMEDIATE) WHEN '1',
	R2O WHEN OTHERS;

	WITH CONTROL(SWITCH_READ_WRITE) SELECT RWSWITCH <= --if SWITCH_READ_WRITE, Read 2 index will be write 1 index
	INSTRUCTION(REGISTER_WRITE_INDEX_1) WHEN '1',
	INSTRUCTION(REGISTER_READ_INDEX_2) WHEN OTHERS;
	
	WITH CONTROL(MEMORY_WRITE_BACK) SELECT REGISTER_WRITEBACK <=
	dDataOut WHEN '1',
	ALU_OUTPUT WHEN OTHERS;

	WITH to_integer(unsigned(INSTRUCTION(REGISTER_WRITE_INDEX_1))) SELECT PC_OVERWRITE <=
	'1' WHEN 31,
	'0' WHEN OTHERS;

	PROCESS (INSTRUCTION(REGISTER_WRITE_INDEX_1),CONTROL(SWITCH_READ_WRITE))
	BEGIN
	IF(to_integer(unsigned(INSTRUCTION(REGISTER_WRITE_INDEX_1))) = 30 AND CONTROL(SWITCH_READ_WRITE) /= '1') THEN
		SP_OVERWRITE <= '1';
	ELSE
		SP_OVERWRITE <= '0';
	END IF;
	END PROCESS;


	PROCESS(CONTROL(POP),CONTROL(PUSH),SP_OUT,ALU_OUTPUT)
		VARIABLE TMP : std_logic_vector(1 downto 0);
	BEGIN
		TMP := CONTROL(POP) & CONTROL(PUSH);
		IF(to_integer(UNSIGNED(TMP)) > 0) THEN
			MEM_ADDRESS <= SP_OUT;
		ELSE
			MEM_ADDRESS <= ALU_OUTPUT;
		END IF;
	END PROCESS;

	WITH to_integer(unsigned(Interrupt_latch & PC_OVERWRITE & CONTROL(JUMP_CONTROL))) SELECT JMP_SELECT <= --Controls branching/changing PC
	'0' WHEN 0,
	'1' WHEN 1,
	Zero_Flag_Latch WHEN 2,
	Carry_Flag_Latch WHEN 3,
	NOT Zero_Flag_Latch WHEN 4,
	'1' WHEN 8, --WHEN PC_OVERWRITE is set
	'1' WHEN 16,
	'0' WHEN OTHERS;

	PROCESS(Interrupt_CPU,Interrupt_latch,CONTROL(MEMORY_TO_PC),dDataOut(9 DOWNTO 0),ALU_OUTPUT(9 DOWNTO 0))
	BEGIN
		IF(Interrupt_CPU = '1' OR Interrupt_latch = '1') THEN
			PC_ALT <= Interrupt_addr;
		ELSIF(CONTROL(MEMORY_TO_PC) = '1') THEN
			PC_ALT <= dDataOut(9 DOWNTO 0);
		ELSE
			PC_ALT <= ALU_OUTPUT(9 DOWNTO 0);
		END IF;
	END PROCESS;

	WITH JMP_SELECT SELECT ADDR <= --Choses instruction to be loaded based on branching
		PC_ALT WHEN '1',
		PC WHEN OTHERS;



	PROCESS  (Interrupt_latch, INSTRUCTION_PRAM)--Changes instruction if interrupt is detected
	BEGIN
		IF(Interrupt_latch = '1') THEN
			INSTRUCTION <= PUSH_PC;
		ELSE
			INSTRUCTION <= INSTRUCTION_PRAM;
		END IF;
	END PROCESS;


	RUN : PROCESS (subClock) --Chose new value of PC based on branching
	BEGIN
		IF (rising_edge(subClock)) THEN --clk
			IF (Interrupt_latch = '1' AND JMP_SELECT /= '1') THEN
				PC <= PC;
			ELSIF (Interrupt_latch = '1' AND JMP_SELECT = '1') THEN
				PC <= PC_ALT;
			ELSIF (JMP_SELECT /= '1') THEN
				PC <= std_logic_vector(unsigned(PC) + 1);
			ELSE
				PC <= std_logic_vector(unsigned(PC_ALT) + 1);
			END IF;
		END IF;
	END PROCESS;

	PROCESS(INSTRUCTION, Interrupt_nest_enable)
	BEGIN
		IF(Interrupt_nest_enable = '0' AND Interrupt_nest_enable_latch = '0') THEN
			Interrupt_enable <= '0';
			Interrupt_nest_enable_latch <= '1';
		ELSIF(INSTRUCTION = POP_PC) THEN
			Interrupt_enable <= '1';
			Interrupt_nest_enable_latch <= '0';
		END IF;
	END PROCESS;

	PROCESS(subClock)
	BEGIN
		IF(rising_edge(subClock)) THEN
			IF(Interrupt_CPU = '1') THEN
				Interrupt_latch <= '1';
				IF(JMP_SELECT = '1') THEN
					PC_INT_TMP <= std_logic_vector(unsigned(PC) - 1);
				ELSE
					PC_INT_TMP <= PC;
				END IF;
			ELSIF(Interrupt_latch = '1') THEN
				Interrupt_latch <= '0';
			END IF;
		END IF;
	END PROCESS;

	--Latches Flags in tempo register, neccesarry due to clock timing
	LATCH : PROCESS (subClock)
	BEGIN
		IF (rising_edge(subClock)) THEN
			Zero_Flag_Latch <= Zero_Flag;
			Overflow_Flag_Latch <= Overflow_Flag;
			Signed_Flag_Latch <= Signed_Flag;
			Parity_Flag_Latch <= Parity_Flag;
			Carry_Flag_Latch <= Carry_Flag;
		END IF;
	END PROCESS;

	PC_REG_IN <= "000000" & std_logic_vector(unsigned(PC) + 1);

--Below controls Clock---

	WITH CONTROL(HALT) SELECT subClock <=
	--PLL_CLOCK_TEMP WHEN '0',
	--DBtn(2) when '0',
	clk when '0',
	'0' WHEN OTHERS;

	WITH PLL_LOCK SELECT PLL_CLOCK_TEMP <=
		PLL_CLOCK WHEN '1',
		'0' WHEN OTHERS;
	PROCESS (PLL_CLOCK)

	BEGIN
		IF (rising_edge(PLL_CLOCK)) THEN
			DIVIDER <= std_logic_vector(unsigned(DIVIDER) + 1);
		END IF;
	END PROCESS;

	btn_inverted <= not btn;

	LED(9) <= Zero_Flag; --Latch not needed
	LED(8) <= Overflow_Flag;
	LED(7) <= Signed_Flag;
	LED(6) <= Parity_Flag;
	LED(5) <= btn_inverted(0);

	LED(0) <= DIVIDER(25);
	LED(1) <= CONTROL(HALT);

END ARCHITECTURE Behavioral;