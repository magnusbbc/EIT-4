Coefs (	std_logic_vector(to_signed(coefs_int(-12),16)), std_logic_vector(to_signed(coefs_int(  -4),16)), std_logic_vector(to_signed(coefs_int(   5),16)), std_logic_vector(to_signed(coefs_int(  17),16)), std_logic_vector(to_signed(coefs_int(  31),16)), std_logic_vector(to_signed(coefs_int(  48),16)), std_logic_vector(to_signed(coefs_int(  65),16)), std_logic_vector(to_signed(coefs_int(  79),16)), std_logic_vector(to_signed(coefs_int(  86, /
       83),16)), std_logic_vector(to_signed(coefs_int(  64),16)), std_logic_vector(to_signed(coefs_int(  26),16)), std_logic_vector(to_signed(coefs_int( -31),16)), std_logic_vector(to_signed(coefs_int(-106),16)), std_logic_vector(to_signed(coefs_int(-194),16)), std_logic_vector(to_signed(coefs_int(-284),16)), std_logic_vector(to_signed(coefs_int(-366),16)), std_logic_vector(to_signed(coefs_int(-424, /
     -442),16)), std_logic_vector(to_signed(coefs_int(-405),16)), std_logic_vector(to_signed(coefs_int(-300),16)), std_logic_vector(to_signed(coefs_int(-120),16)), std_logic_vector(to_signed(coefs_int( 139),16)), std_logic_vector(to_signed(coefs_int( 470),16)), std_logic_vector(to_signed(coefs_int( 862),16)), std_logic_vector(to_signed(coefs_int(1295),16)), std_logic_vector(to_signed(coefs_int(1744, /
     2182),16)), std_logic_vector(to_signed(coefs_int(2578),16)), std_logic_vector(to_signed(coefs_int(2904),16)), std_logic_vector(to_signed(coefs_int(3137),16)), std_logic_vector(to_signed(coefs_int(3256),16)), std_logic_vector(to_signed(coefs_int(3257),16)), std_logic_vector(to_signed(coefs_int(3137),16)), std_logic_vector(to_signed(coefs_int(2904),16)), std_logic_vector(to_signed(coefs_int(2578, /
     2182),16)), std_logic_vector(to_signed(coefs_int(1744),16)), std_logic_vector(to_signed(coefs_int(1295),16)), std_logic_vector(to_signed(coefs_int( 862),16)), std_logic_vector(to_signed(coefs_int( 470),16)), std_logic_vector(to_signed(coefs_int( 139),16)), std_logic_vector(to_signed(coefs_int(-120),16)), std_logic_vector(to_signed(coefs_int(-300),16)), std_logic_vector(to_signed(coefs_int(-405, /
     -442),16)), std_logic_vector(to_signed(coefs_int(-424),16)), std_logic_vector(to_signed(coefs_int(-366),16)), std_logic_vector(to_signed(coefs_int(-284),16)), std_logic_vector(to_signed(coefs_int(-194),16)), std_logic_vector(to_signed(coefs_int(-106),16)), std_logic_vector(to_signed(coefs_int( -31),16)), std_logic_vector(to_signed(coefs_int(  26),16)), std_logic_vector(to_signed(coefs_int(  64, / 
       83),16)), std_logic_vector(to_signed(coefs_int(  86),16)), std_logic_vector(to_signed(coefs_int(  79),16)), std_logic_vector(to_signed(coefs_int(  65),16)), std_logic_vector(to_signed(coefs_int(  48),16)), std_logic_vector(to_signed(coefs_int(  31),16)), std_logic_vector(to_signed(coefs_int(  17),16)), std_logic_vector(to_signed(coefs_int(   5),16)), std_logic_vector(to_signed(coefs_int(  -4, /
      -12); /