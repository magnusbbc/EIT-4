Multiplier_1_inst : Multiplier_1 PORT MAP (
		dataa	 => dataa_sig,
		datab	 => datab_sig,
		result	 => result_sig
	);
